��(4      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �min_impurity_split�N�class_weight�N�	ccp_alpha�G        �_sklearn_version��0.24.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hNhG        �n_features_in_�K�n_features_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h-�dtype����i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��h6�f8�����R�(Kh:NNNJ����J����K t�b�C              �?�t�bh>h*�scalar���h9C       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hK�
node_count�K�nodes�h,h/K ��h1��R�(KK��h6�V56�����R�(K�|�N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hkh9K ��hlh9K��hmh9K��hnhJK��hohJK ��hph9K(��hqhJK0��uK8KKt�b�BH                              @�q�q�?(            �O@������������������������       �                     A@                           �?�c�Α�?             =@                          ph@��S���?             .@                          �5@�<ݚ�?             "@������������������������       �                     �?                            @      �?              @       	                 ���f@���Q��?             @������������������������       �                     �?
                          �g@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             ,@�t�b�values�h,h/K ��h1��R�(KKKK��hJ�C�      E@      5@      A@               @      5@       @      @       @      @              �?       @      @       @      @      �?              �?      @              @      �?                      @      @                      ,@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�BH                              @���h%��?*            �O@������������������������       �                    �C@                        ���e@r�q��?             8@������������������������       �                      @       
                 ���f@�C��2(�?             6@                          �5@      �?             @������������������������       �                      @       	                    H@      �?              @������������������������       �                     �?������������������������       �                     �?                            @�X�<ݺ?             2@                          �g@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             *@�t�bh~h,h/K ��h1��R�(KKKK��hJ�C�     �E@      4@     �C@              @      4@       @               @      4@      �?      @               @      �?      �?      �?                      �?      �?      1@      �?      @              @      �?                      *@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK	hbh,h/K ��h1��R�(KK	��hi�B�                              @�ՙ/�?'            �O@������������������������       �                    �@@                            @z�G�z�?             >@                          �g@���Q��?
             .@                        ���f@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     @������������������������       �        	             .@�t�bh~h,h/K ��h1��R�(KK	KK��hJ�C�     �C@      8@     �@@              @      8@      @      "@      �?      "@      �?                      "@      @                      .@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaK	hbh,h/K ��h1��R�(KK	��hi�B�                              @b����?&            �O@                            @�:�^���?            �F@������������������������       �                    �A@                          �g@���Q��?             $@                          �@@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     2@�t�bh~h,h/K ��h1��R�(KK	KK��hJ�C�     �D@      6@     �D@      @     �A@              @      @       @      @       @                      @      @                      2@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�Bh                              @�ՙ/�?+            �O@������������������������       �                    �@@       
                     @z�G�z�?             >@       	                 0E�D@      �?             (@                          �g@      �?              @                        ���f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     2@�t�bh~h,h/K ��h1��R�(KKKK��hJ�C�     �C@      8@     �@@              @      8@      @      @      @       @      �?       @      �?                       @      @                      @              2@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�B�                            0f@��~R���?)            �O@                           �?���7�?             6@������������������������       �                     4@                          �I@      �?              @������������������������       �                     �?������������������������       �                     �?       
                   �g@D^��#��?            �D@       	                     @�q�q�?             8@������������������������       �                     ,@������������������������       �                     $@                        0E~B@�t����?             1@                            @8�Z$���?             *@������������������������       �                      @������������������������       �                     &@                           @      �?             @������������������������       �                     @������������������������       �                     �?�t�bh~h,h/K ��h1��R�(KKKK��hJ�B        D@      7@      5@      �?      4@              �?      �?      �?                      �?      3@      6@      ,@      $@      ,@                      $@      @      (@       @      &@       @                      &@      @      �?      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�B�                            �d@�ՙ/�?&            �O@������������������������       �        	             ,@                            @�`���?            �H@������������������������       �                     6@                            @�����H�?             ;@                           h@      �?              @       
                 ���f@r�q��?             @       	                    H@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     3@�t�bh~h,h/K ��h1��R�(KKKK��hJ�C�     �C@      8@      ,@              9@      8@      6@              @      8@      @      @      �?      @      �?      @      �?                      @               @       @                      3@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�Bh                              @��~R���?*            �O@������������������������       �                     @@       
                 0E�D@r֛w���?             ?@       	                     @���Q��?             4@                          �g@�n_Y�K�?             *@                        ���f@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     &@�t�bh~h,h/K ��h1��R�(KKKK��hJ�C�      D@      7@      @@               @      7@       @      (@       @      @      �?      @      �?                      @      @                      @              &@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�BH                            0f@p�EG/��?,            �O@                            @�C��2(�?             6@������������������������       �                     4@������������������������       �                      @                            @�>$�*��?            �D@                           @ �o_��?             9@                            @؇���X�?             5@������������������������       �                     $@	                          �g@���!pc�?             &@
                        ���f@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     0@�t�bh~h,h/K ��h1��R�(KKKK��hJ�C�      C@      9@      4@       @      4@                       @      2@      7@      2@      @      2@      @      $@               @      @      @      @      @                      @      @                      @              0@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhNhG        h'Kh&Kh(Kh)h,h/K ��h1��R�(KK��hJ�C              �?�t�bh>hOh9C       ���R�hSKhThWKh,h/K ��h1��R�(KK��h9�C       �t�bK��R�}�(hKhaKhbh,h/K ��h1��R�(KK��hi�Bh                              @������?%            �O@������������������������       �                     :@       
                    �?$G$n��?            �B@       	                     @���N8�?             5@                          �g@      �?              @                          0f@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     *@������������������������       �        	             0@�t�bh~h,h/K ��h1��R�(KKKK��hJ�C�      ?@      @@      :@              @      @@      @      0@      @      @       @      @       @                      @      @                      *@              0@�t�bubhhubehhub.